/* The 32x32-bit S-Box S1
* Input: a 32-bit input.
* Output: a 32-bit output of S1 box.
*/
module S1(
  input  [31:0] w,
  input clk,
  output [31:0] s1_out
);
  
  reg [7:0] SR [0:255];
  reg [31:0] r0, r1, r2, r3;
  
  reg [7:0] srw0, srw1, srw2, srw3;
  wire [7:0] mulx_out0, mulx_out1, mulx_out2, mulx_out3;

  MULx MULx_0(.V(srw0), .c(8'h1b),.clk(clk), .mulx_out(mulx_out0)); 
  MULx MULx_1(.V(srw1), .c(8'h1b),.clk(clk), .mulx_out(mulx_out1));
  MULx MULx_2(.V(srw2), .c(8'h1b),.clk(clk), .mulx_out(mulx_out2));
  MULx MULx_3(.V(srw3), .c(8'h1b),.clk(clk), .mulx_out(mulx_out3));
 
  always @(*) begin

    // Initializing SR 
    SR[0]   = 8'h63;
    SR[1]   = 8'h7C;
    SR[2]   = 8'h77;
    SR[3]   = 8'h7B;
    SR[4]   = 8'hF2;
    SR[5]   = 8'h6B;
    SR[6]   = 8'h6F;
    SR[7]   = 8'hC5;
    SR[8]   = 8'h30;
    SR[9]   = 8'h01;
    SR[10]  = 8'h67;
    SR[11]  = 8'h2B;
    SR[12]  = 8'hFE;
    SR[13]  = 8'hD7;
    SR[14]  = 8'hAB;
    SR[15]  = 8'h76;
    SR[16]  = 8'hCA;
    SR[17]  = 8'h82;
    SR[18]  = 8'hC9;
    SR[19]  = 8'h7D;
    SR[20]  = 8'hFA;
    SR[21]  = 8'h59;
    SR[22]  = 8'h47;
    SR[23]  = 8'hF0;
    SR[24]  = 8'hAD;
    SR[25]  = 8'hD4;
    SR[26]  = 8'hA2;
    SR[27]  = 8'hAF;
    SR[28]  = 8'h9C;
    SR[29]  = 8'hA4;
    SR[30]  = 8'h72;
    SR[31]  = 8'hC0;
    SR[32]  = 8'hB7;
    SR[33]  = 8'hFD;
    SR[34]  = 8'h93;
    SR[35]  = 8'h26;
    SR[36]  = 8'h36;
    SR[37]  = 8'h3F;
    SR[38]  = 8'hF7;
    SR[39]  = 8'hCC;
    SR[40]  = 8'h34;
    SR[41]  = 8'hA5;
    SR[42]  = 8'hE5;
    SR[43]  = 8'hF1;
    SR[44]  = 8'h71;
    SR[45]  = 8'hD8;
    SR[46]  = 8'h31;
    SR[47]  = 8'h15;
    SR[48]  = 8'h04;
    SR[49]  = 8'hC7;
    SR[50]  = 8'h23;
    SR[51]  = 8'hC3;
    SR[52]  = 8'h18;
    SR[53]  = 8'h96;
    SR[54]  = 8'h05;
    SR[55]  = 8'h9A;
    SR[56]  = 8'h07;
    SR[57]  = 8'h12;
    SR[58]  = 8'h80;
    SR[59]  = 8'hE2;
    SR[60]  = 8'hEB;
    SR[61]  = 8'h27;
    SR[62]  = 8'hB2;
    SR[63]  = 8'h75;
    SR[64]  = 8'h09;
    SR[65]  = 8'h83;
    SR[66]  = 8'h2C;
    SR[67]  = 8'h1A;
    SR[68]  = 8'h1B;
    SR[69]  = 8'h6E;
    SR[70]  = 8'h5A;
    SR[71]  = 8'hA0;
    SR[72]  = 8'h52;
    SR[73]  = 8'h3B;
    SR[74]  = 8'hD6;
    SR[75]  = 8'hB3;
    SR[76]  = 8'h29;
    SR[77]  = 8'hE3;
    SR[78]  = 8'h2F;
    SR[79]  = 8'h84;
    SR[80]  = 8'h53;
    SR[81]  = 8'hD1;
    SR[82]  = 8'h00;
    SR[83]  = 8'hED;
    SR[84]  = 8'h20;
    SR[85]  = 8'hFC;
    SR[86]  = 8'hB1;
    SR[87]  = 8'h5B;
    SR[88]  = 8'h6A;
    SR[89]  = 8'hCB;
    SR[90]  = 8'hBE;
    SR[91]  = 8'h39;
    SR[92]  = 8'h4A;
    SR[93]  = 8'h4C;
    SR[94]  = 8'h58;
    SR[95]  = 8'hCF;
    SR[96]  = 8'hD0;
    SR[97]  = 8'hEF;
    SR[98]  = 8'hAA;
    SR[99]  = 8'hFB;
    SR[100] = 8'h43;
    SR[101] = 8'h4D;
    SR[102] = 8'h33;
    SR[103] = 8'h85;
    SR[104] = 8'h45;
    SR[105] = 8'hF9;
    SR[106] = 8'h02;
    SR[107] = 8'h7F;
    SR[108] = 8'h50;
    SR[109] = 8'h3C;
    SR[110] = 8'h9F;
    SR[111] = 8'hA8;
    SR[112] = 8'h51;
    SR[113] = 8'hA3;
    SR[114] = 8'h40;
    SR[115] = 8'h8F;
    SR[116] = 8'h92;
    SR[117] = 8'h9D;
    SR[118] = 8'h38;
    SR[119] = 8'hF5;
    SR[120] = 8'hBC;
    SR[121] = 8'hB6;
    SR[122] = 8'hDA;
    SR[123] = 8'h21;
    SR[124] = 8'h10;
    SR[125] = 8'hFF;
    SR[126] = 8'hF3;
    SR[127] = 8'hD2;
    SR[128] = 8'hCD;
    SR[129] = 8'h0C;
    SR[130] = 8'h13;
    SR[131] = 8'hEC;
    SR[132] = 8'h5F;
    SR[133] = 8'h97;
    SR[134] = 8'h44;
    SR[135] = 8'h17;
    SR[136] = 8'hC4;
    SR[137] = 8'hA7;
    SR[138] = 8'h7E;
    SR[139] = 8'h3D;
    SR[140] = 8'h64;
    SR[141] = 8'h5D;
    SR[142] = 8'h19;
    SR[143] = 8'h73;
    SR[144] = 8'h60;
    SR[145] = 8'h81;
    SR[146] = 8'h4F;
    SR[147] = 8'hDC;
    SR[148] = 8'h22;
    SR[149] = 8'h2A;
    SR[150] = 8'h90;
    SR[151] = 8'h88;
    SR[152] = 8'h46;
    SR[153] = 8'hEE;
    SR[154] = 8'hB8;
    SR[155] = 8'h14;
    SR[156] = 8'hDE;
    SR[157] = 8'h5E;
    SR[158] = 8'h0B;
    SR[159] = 8'hDB;
    SR[160] = 8'hE0;
    SR[161] = 8'h32;
    SR[162] = 8'h3A;
    SR[163] = 8'h0A;
    SR[164] = 8'h49;
    SR[165] = 8'h06;
    SR[166] = 8'h24;
    SR[167] = 8'h5C;
    SR[168] = 8'hC2;
    SR[169] = 8'hD3;
    SR[170] = 8'hAC;
    SR[171] = 8'h62;
    SR[172] = 8'h91;
    SR[173] = 8'h95;
    SR[174] = 8'hE4;
    SR[175] = 8'h79;
    SR[176] = 8'hE7;
    SR[177] = 8'hC8;
    SR[178] = 8'h37;
    SR[179] = 8'h6D;
    SR[180] = 8'h8D;
    SR[181] = 8'hD5;
    SR[182] = 8'h4E;
    SR[183] = 8'hA9;
    SR[184] = 8'h6C;
    SR[185] = 8'h56;
    SR[186] = 8'hF4;
    SR[187] = 8'hEA;
    SR[188] = 8'h65;
    SR[189] = 8'h7A;
    SR[190] = 8'hAE;
    SR[191] = 8'h08;
    SR[192] = 8'hBA;
    SR[193] = 8'h78;
    SR[194] = 8'h25;
    SR[195] = 8'h2E;
    SR[196] = 8'h1C;
    SR[197] = 8'hA6;
    SR[198] = 8'hB4;
    SR[199] = 8'hC6;
    SR[200] = 8'hE8;
    SR[201] = 8'hDD;
    SR[202] = 8'h74;
    SR[203] = 8'h1F;
    SR[204] = 8'h4B;
    SR[205] = 8'hBD;
    SR[206] = 8'h8B;
    SR[207] = 8'h8A;
    SR[208] = 8'h70;
    SR[209] = 8'h3E;
    SR[210] = 8'hB5;
    SR[211] = 8'h66;
    SR[212] = 8'h48;
    SR[213] = 8'h03;
    SR[214] = 8'hF6;
    SR[215] = 8'h0E;
    SR[216] = 8'h61;
    SR[217] = 8'h35;
    SR[218] = 8'h57;
    SR[219] = 8'hB9;
    SR[220] = 8'h86;
    SR[221] = 8'hC1;
    SR[222] = 8'h1D;
    SR[223] = 8'h9E;
    SR[224] = 8'hE1;
    SR[225] = 8'hF8;
    SR[226] = 8'h98;
    SR[227] = 8'h11;
    SR[228] = 8'h69;
    SR[229] = 8'hD9;
    SR[230] = 8'h8E;
    SR[231] = 8'h94;
    SR[232] = 8'h9B;
    SR[233] = 8'h1E;
    SR[234] = 8'h87;
    SR[235] = 8'hE9;
    SR[236] = 8'hCE;
    SR[237] = 8'h55;
    SR[238] = 8'h28;
    SR[239] = 8'hDF;
    SR[240] = 8'h8C;
    SR[241] = 8'hA1;
    SR[242] = 8'h89;
    SR[243] = 8'h0D;
    SR[244] = 8'hBF;
    SR[245] = 8'hE6;
    SR[246] = 8'h42;
    SR[247] = 8'h68;
    SR[248] = 8'h41;
    SR[249] = 8'h99;
    SR[250] = 8'h2D;
    SR[251] = 8'h0F;
    SR[252] = 8'hB0;
    SR[253] = 8'h54;
    SR[254] = 8'hBB;
    SR[255] = 8'h16;

    
    srw0 = SR[ (w >> 24) & 8'hff ];
    srw1 = SR[ (w >> 16) & 8'hff ];
    srw2 = SR[ (w >> 8) & 8'hff] ;
    srw3 = SR[ w & 8'hff ];
    
    
    r0 = ( ( mulx_out0 ) ^ srw1 ) ^ srw2 ^ ( ( mulx_out3) ) ^ srw3 ;
    r1 = ( ( ( mulx_out0 ) ^ srw0 ) ^ ( mulx_out1 ) ) ^ srw2 ^ srw3;
    r2 = ( srw0 ^ ( ( mulx_out1 ) ^ srw1 ) ^ ( mulx_out2 ) ) ^ srw3;
    r3 = ( srw0 ^ srw1 ) ^ ( ( mulx_out2 ) ^ srw2 ) ^ ( mulx_out3 );

  end
  assign s1_out = ( ( r0 << 24 ) | ( r1 << 16 ) | ( r2 << 8 ) | r3 );
  
endmodule