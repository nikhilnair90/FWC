/* The 32x32-bit S-Box S2
* Input: a 32-bit input.
* Output: a 32-bit output of S2 box.
*/
module S2(
  input  [31:0] w,
  input clk,
  output [31:0] s2_out
);
    
  reg [7:0] SQ [0:255];
  reg [31:0] r0, r1, r2, r3;
  
  reg [7:0] sqw0, sqw1, sqw2, sqw3;
  wire [7:0] mulx_out4, mulx_out5, mulx_out6, mulx_out7;

  MULx MULx_0(.V(sqw0), .c(8'h69),.clk(clk), .mulx_out(mulx_out4)); 
  MULx MULx_1(.V(sqw1), .c(8'h69),.clk(clk), .mulx_out(mulx_out5));
  MULx MULx_2(.V(sqw2), .c(8'h69),.clk(clk), .mulx_out(mulx_out6));
  MULx MULx_3(.V(sqw3), .c(8'h69),.clk(clk), .mulx_out(mulx_out7));
 
  always @(*) begin

     //Initializing SQ
    SQ[0]   = 8'h25;
    SQ[1]   = 8'h24;
    SQ[2]   = 8'h73;
    SQ[3]   = 8'h67;
    SQ[4]   = 8'hD7;
    SQ[5]   = 8'hAE;
    SQ[6]   = 8'h5C;
    SQ[7]   = 8'h30;
    SQ[8]   = 8'hA4;
    SQ[9]   = 8'hEE;
    SQ[10]  = 8'h6E;
    SQ[11]  = 8'hCB;
    SQ[12]  = 8'h7D;
    SQ[13]  = 8'hB5;
    SQ[14]  = 8'h82;
    SQ[15]  = 8'hDB;
    SQ[16]  = 8'hE4;
    SQ[17]  = 8'h8E;
    SQ[18]  = 8'h48;
    SQ[19]  = 8'h49;
    SQ[20]  = 8'h4F;
    SQ[21]  = 8'h5D;
    SQ[22]  = 8'h6A;
    SQ[23]  = 8'h78;
    SQ[24]  = 8'h70;
    SQ[25]  = 8'h88;
    SQ[26]  = 8'hE8;
    SQ[27]  = 8'h5F;
    SQ[28]  = 8'h5E;
    SQ[29]  = 8'h84;
    SQ[30]  = 8'h65;
    SQ[31]  = 8'hE2;
    SQ[32]  = 8'hD8;
    SQ[33]  = 8'hE9;
    SQ[34]  = 8'hCC;
    SQ[35]  = 8'hED;
    SQ[36]  = 8'h40;
    SQ[37]  = 8'h2F;
    SQ[38]  = 8'h11;
    SQ[39]  = 8'h28;
    SQ[40]  = 8'h57;
    SQ[41]  = 8'hD2;
    SQ[42]  = 8'hAC;
    SQ[43]  = 8'hE3;
    SQ[44]  = 8'h4A;
    SQ[45]  = 8'h15;
    SQ[46]  = 8'h1B;
    SQ[47]  = 8'hB9;
    SQ[48]  = 8'hB2;
    SQ[49]  = 8'h80;
    SQ[50]  = 8'h85;
    SQ[51]  = 8'hA6;
    SQ[52]  = 8'h2E;
    SQ[53]  = 8'h02;
    SQ[54]  = 8'h47;
    SQ[55]  = 8'h29;
    SQ[56]  = 8'h07;
    SQ[57]  = 8'h4B;
    SQ[58]  = 8'h0E;
    SQ[59]  = 8'hC1;
    SQ[60]  = 8'h51;
    SQ[61]  = 8'hAA;
    SQ[62]  = 8'h89;
    SQ[63]  = 8'hD4;
    SQ[64]  = 8'hCA;
    SQ[65]  = 8'h01;
    SQ[66]  = 8'h46;
    SQ[67]  = 8'hB3;
    SQ[68]  = 8'hEF;
    SQ[69]  = 8'hDD;
    SQ[70]  = 8'h44;
    SQ[71]  = 8'h7B;
    SQ[72]  = 8'hC2;
    SQ[73]  = 8'h7F;
    SQ[74]  = 8'hBE;
    SQ[75]  = 8'hC3;
    SQ[76]  = 8'h9F;
    SQ[77]  = 8'h20;
    SQ[78]  = 8'h4C;
    SQ[79]  = 8'h64;
    SQ[80]  = 8'h83;
    SQ[81]  = 8'hA2;
    SQ[82]  = 8'h68;
    SQ[83]  = 8'h42;
    SQ[84]  = 8'h13;
    SQ[85]  = 8'hB4;
    SQ[86]  = 8'h41;
    SQ[87]  = 8'hCD;
    SQ[88]  = 8'hBA;
    SQ[89]  = 8'hC6;
    SQ[90]  = 8'hBB;
    SQ[91]  = 8'h6D;
    SQ[92]  = 8'h4D;
    SQ[93]  = 8'h71;
    SQ[94]  = 8'h21;
    SQ[95]  = 8'hF4;
    SQ[96]  = 8'h8D;
    SQ[97]  = 8'hB0;
    SQ[98]  = 8'hE5;
    SQ[99]  = 8'h93;
    SQ[100] = 8'hFE;
    SQ[101] = 8'h8F;
    SQ[102] = 8'hE6;
    SQ[103] = 8'hCF;
    SQ[104] = 8'h43;
    SQ[105] = 8'h45;
    SQ[106] = 8'h31;
    SQ[107] = 8'h22;
    SQ[108] = 8'h37;
    SQ[109] = 8'h36;
    SQ[110] = 8'h96;
    SQ[111] = 8'hFA;
    SQ[112] = 8'hBC;
    SQ[113] = 8'h0F;
    SQ[114] = 8'h08;
    SQ[115] = 8'h52;
    SQ[116] = 8'h1D;
    SQ[117] = 8'h55;
    SQ[118] = 8'h1A;
    SQ[119] = 8'hC5;
    SQ[120] = 8'h4E;
    SQ[121] = 8'h23;
    SQ[122] = 8'h69;
    SQ[123] = 8'h7A;
    SQ[124] = 8'h92;
    SQ[125] = 8'hFF;
    SQ[126] = 8'h5B;
    SQ[127] = 8'h5A;
    SQ[128] = 8'hEB;
    SQ[129] = 8'h9A;
    SQ[130] = 8'h1C;
    SQ[131] = 8'hA9;
    SQ[132] = 8'hD1;
    SQ[133] = 8'h7E;
    SQ[134] = 8'h0D;
    SQ[135] = 8'hFC;
    SQ[136] = 8'h50;
    SQ[137] = 8'h8A;
    SQ[138] = 8'hB6;
    SQ[139] = 8'h62;
    SQ[140] = 8'hF5;
    SQ[141] = 8'h0A;
    SQ[142] = 8'hF8;
    SQ[143] = 8'hDC;
    SQ[144] = 8'h03;
    SQ[145] = 8'h3C;
    SQ[146] = 8'h0C;
    SQ[147] = 8'h39;
    SQ[148] = 8'hF1;
    SQ[149] = 8'hB8;
    SQ[150] = 8'hF3;
    SQ[151] = 8'h3D;
    SQ[152] = 8'hF2;
    SQ[153] = 8'hD5;
    SQ[154] = 8'h97;
    SQ[155] = 8'h66;
    SQ[156] = 8'h81;
    SQ[157] = 8'h32;
    SQ[158] = 8'hA0;
    SQ[159] = 8'h00;
    SQ[160] = 8'h06;
    SQ[161] = 8'hCE;
    SQ[162] = 8'hF6;
    SQ[163] = 8'hEA;
    SQ[164] = 8'hB7;
    SQ[165] = 8'h17;
    SQ[166] = 8'hF7;
    SQ[167] = 8'h8C;
    SQ[168] = 8'h79;
    SQ[169] = 8'hD6;
    SQ[170] = 8'hA7;
    SQ[171] = 8'hBF;
    SQ[172] = 8'h8B;
    SQ[173] = 8'h3F;
    SQ[174] = 8'h1F;
    SQ[175] = 8'h53;
    SQ[176] = 8'h63;
    SQ[177] = 8'h75;
    SQ[178] = 8'h35;
    SQ[179] = 8'h2C;
    SQ[180] = 8'h60;
    SQ[181] = 8'hFD;
    SQ[182] = 8'h27;
    SQ[183] = 8'hD3;
    SQ[184] = 8'h94;
    SQ[185] = 8'hA5;
    SQ[186] = 8'h7C;
    SQ[187] = 8'hA1;
    SQ[188] = 8'h05;
    SQ[189] = 8'h58;
    SQ[190] = 8'h2D;
    SQ[191] = 8'hBD;
    SQ[192] = 8'hD9;
    SQ[193] = 8'hC7;
    SQ[194] = 8'hAF;
    SQ[195] = 8'h6B;
    SQ[196] = 8'h54;
    SQ[197] = 8'h0B;
    SQ[198] = 8'hE0;
    SQ[199] = 8'h38;
    SQ[200] = 8'h04;
    SQ[201] = 8'hC8;
    SQ[202] = 8'h9D;
    SQ[203] = 8'hE7;
    SQ[204] = 8'h14;
    SQ[205] = 8'hB1;
    SQ[206] = 8'h87;
    SQ[207] = 8'h9C;
    SQ[208] = 8'hDF;
    SQ[209] = 8'h6F;
    SQ[210] = 8'hF9;
    SQ[211] = 8'hDA;
    SQ[212] = 8'h2A;
    SQ[213] = 8'hC4;
    SQ[214] = 8'h59;
    SQ[215] = 8'h16;
    SQ[216] = 8'h74;
    SQ[217] = 8'h91;
    SQ[218] = 8'hAB;
    SQ[219] = 8'h26;
    SQ[220] = 8'h61;
    SQ[221] = 8'h76;
    SQ[222] = 8'h34;
    SQ[223] = 8'h2B;
    SQ[224] = 8'hAD;
    SQ[225] = 8'h99;
    SQ[226] = 8'hFB;
    SQ[227] = 8'h72;
    SQ[228] = 8'hEC;
    SQ[229] = 8'h33;
    SQ[230] = 8'h12;
    SQ[231] = 8'hDE;
    SQ[232] = 8'h98;
    SQ[233] = 8'h3B;
    SQ[234] = 8'hC0;
    SQ[235] = 8'h9B;
    SQ[236] = 8'h3E;
    SQ[237] = 8'h18;
    SQ[238] = 8'h10;
    SQ[239] = 8'h3A;
    SQ[240] = 8'h56;
    SQ[241] = 8'hE1;
    SQ[242] = 8'h77;
    SQ[243] = 8'hC9;
    SQ[244] = 8'h1E;
    SQ[245] = 8'h9E;
    SQ[246] = 8'h95;
    SQ[247] = 8'hA3;
    SQ[248] = 8'h90;
    SQ[249] = 8'h19;
    SQ[250] = 8'hA8;
    SQ[251] = 8'h6C;
    SQ[252] = 8'h09;
    SQ[253] = 8'hD0;
    SQ[254] = 8'hF0;
    SQ[255] = 8'h86;


    
    sqw0 = SQ[ (w >> 24) & 8'hff ];
    sqw1 = SQ[ (w >> 16) & 8'hff ];
    sqw2 = SQ[ (w >> 8) & 8'hff] ;
    sqw3 = SQ[ w & 8'hff ];
    
    r0 = ( ( mulx_out4 ) ^ sqw1 ) ^ sqw2 ^ ( ( mulx_out7) ) ^ sqw3 ;
    r1 = ( ( ( mulx_out4 ) ^ sqw0 ) ^ ( mulx_out5 ) ) ^ sqw2 ^ sqw3;
    r2 = ( sqw0 ^ ( ( mulx_out5 ) ^ sqw1 ) ^ ( mulx_out6 ) ) ^ sqw3;
    r3 = ( sqw0 ^ sqw1 ) ^ ( ( mulx_out6 ) ^ sqw2 ) ^ ( mulx_out7 );
    
    
  end
  assign s2_out = ( ( r0 << 24 ) | ( r1 << 16 ) | ( r2 << 8 ) | r3 );
  
endmodule